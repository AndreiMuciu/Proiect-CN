library verilog;
use verilog.vl_types.all;
entity CSkA_tb is
    generic(
        N               : integer := 32
    );
end CSkA_tb;
